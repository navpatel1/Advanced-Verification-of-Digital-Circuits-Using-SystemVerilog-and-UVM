// module mux
//   (
//     input [3:0] a,b,c,d, ////input data port have size of 4-bit
//     input [1:0] sel,     ////control port have size of 2-bit
//     output reg [3:0] y 
//   );
  
//   always@(*)
//     begin
//       case(sel)
//         2'b00: y = a;
//         2'b01: y = b;
//         2'b10: y = c;
//         2'b11: y = d;
//       endcase
//     end
  
  
// endmodule
// Questions for this assignment
// Design UVM testbench to perform verification of 4:1 Mux. Design code of 4:1 Mux is added in the Instruction tab.


